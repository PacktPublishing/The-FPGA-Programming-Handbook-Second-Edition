../../../CH6/SystemVerilog/tb/adt7420_mdl.sv