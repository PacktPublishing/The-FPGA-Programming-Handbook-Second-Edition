../../../CH6/SystemVerilog/tb/tb_temp.sv